////////////////////////////////////////////////////////////////
// Copyright (c) 2019 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
////////////////////////////////////////////////////////////////
//Description:
//Author:  wxxiao
//History: v1.0
////////////////////////////////////////////////////////////////
`timescale 1ns/1ps
module ips2l_ddrphy_ppll_v1_0 #(
parameter  real CLKIN_FREQ =  50.0,
parameter  BANDWIDTH      = "OPTIMIZED",
parameter  CLKOUT4_SYN_EN = "FLASE",
parameter  INTERNAL_FB    = "CLKOUTF",
parameter  IDIV           =  2,
parameter  FDIV           =  64,
parameter  ODIVPHY        =  4      //8'd2:800  8'd4:400
)(
input   clk_in0,
input   pll_rst,
input   clkoutphy_gate,
output  clkout0,
output  clkout0n,
output  clkoutphy,
output  clkoutphyn,
output  pll_lock
);

parameter   ODIV0   =  16;    //100
parameter   ODIV1   =  2;
parameter   ODIV2   =  4;
parameter   ODIV3   =  8;
parameter   ODIV4   =  FDIV/IDIV;

GTP_PPLL #(
   .CLKIN_FREQ         (CLKIN_FREQ),   
   .LOCK_MODE          (1'b0   ),      
   .STATIC_RATIOI      (IDIV   ),      
   .STATIC_RATIOM      (1      ),      
   .STATIC_RATIO0      (ODIV0  ),      
   .STATIC_RATIO1      (ODIV1  ),      
   .STATIC_RATIO2      (ODIV2  ),      
   .STATIC_RATIO3      (ODIV3  ),      
   .STATIC_RATIO4      (ODIV4  ),      
   .STATIC_RATIOPHY    (ODIVPHY),      
   .STATIC_RATIOF      (FDIV   ),      
   .STATIC_DUTY0       (ODIV0  ),      
   .STATIC_DUTY1       (ODIV1  ),      
   .STATIC_DUTY2       (ODIV2  ),      
   .STATIC_DUTY3       (ODIV3  ),      
   .STATIC_DUTY4       (ODIV4  ),      
   .STATIC_DUTYPHY     (ODIVPHY),      
   .STATIC_DUTYF       (FDIV   ),      
   .STATIC_PHASE0      (0),            
   .STATIC_PHASE1      (0),            
   .STATIC_PHASE2      (0),            
   .STATIC_PHASE3      (0),            
   .STATIC_PHASE4      (0),            
   .STATIC_PHASEPHY    (0),            
   .STATIC_PHASEF      (0),            
   .STATIC_CPHASE0     (0),            
   .STATIC_CPHASE1     (0),            
   .STATIC_CPHASE2     (0),            
   .STATIC_CPHASE3     (0),            
   .STATIC_CPHASE4     (0),            
   .STATIC_CPHASEPHY   (0),            
   .STATIC_CPHASEF     (0),            
   .CLKOUT0_SYN_EN     ("FALSE"),      
   .CLKOUT1_SYN_EN     ("FALSE"),      
   .CLKOUT2_SYN_EN     ("FALSE"),      
   .CLKOUT3_SYN_EN     ("FALSE"),      
   .CLKOUT4_SYN_EN     (CLKOUT4_SYN_EN),
   .CLKOUTPHY_SYN_EN   ("TRUE"),       
   .CLKOUTF_SYN_EN     ("FALSE"),      
   .INTERNAL_FB        (INTERNAL_FB) ,
   .EXTERNAL_FB        ("DISABLE"),    
   .BANDWIDTH          (BANDWIDTH)   
    )u_ppll(
   .CLKOUT0          (clkout0   ),               
   .CLKOUT0N         (clkout0n  ),
   .CLKOUT1          (),
   .CLKOUT1N         (),
   .CLKOUT2          (),
   .CLKOUT2N         (),
   .CLKOUT3          (),
   .CLKOUT3N         (),
   .CLKOUT4          (),
   .CLKOUTPHY        (clkoutphy),
   .CLKOUTPHYN       (clkoutphyn),
   .CLKOUTF          (),
   .CLKOUTFN         (),
   .LOCK             (pll_lock),
   .APB_RDATA        (),
   .APB_READY        (),
   .CLKIN1           (clk_in0),
   .CLKIN2           (1'b0),
   .CLKFB            (1'b0),
   .CLKIN_SEL        (1'b0),
   .CLKOUT0_SYN      (1'b0),
   .CLKOUT1_SYN      (1'b0),
   .CLKOUT2_SYN      (1'b0),
   .CLKOUT3_SYN      (1'b0),
   .CLKOUT4_SYN      (1'b0),
   .CLKOUTPHY_SYN    (clkoutphy_gate),
   .CLKOUTF_SYN      (1'b0),
   .PLL_PWD          (1'b0),
   .RST              (pll_rst),
   .APB_CLK          (1'b0),
   .APB_RST_N        (1'b0),
   .APB_ADDR         (5'd0),
   .APB_SEL          (1'b0),
   .APB_EN           (1'b0),
   .APB_WRITE        (1'b0),
   .APB_WDATA        (16'd0)
    );

//   PPLL u_ppll( 
//     .SC_ALDO_LOAD_CTRL                 (1'b0),
//     .SC_ALDO_LPF_ADJ                   (2'b00),
//     .SC_ALDO_TEST                      (2'b11),
//     .SC_ALDO_TEST_EN                   (1'b0),
//     .SC_ALDO_VREF_ADJ                  (3'b000),
//     .SC_ALDO_VREF_SEL                  (4'b0000),
//     .SC_CLKFBOUT_GATE_EN               (1'b0),
//     .SC_CLKINORFB_DLYSEL               (2'b00),
//     .SC_CLKINORFB_DLYSET               (6'd0),
//     .SC_CLKIN_STASEL                   (1'b0),
//     .SC_CLKOUT0_GATE_EN                (1'b0),
//     .SC_CLKOUT1_GATE_EN                (1'b0),
//     .SC_CLKOUT2_GATE_EN                (1'b0),
//     .SC_CLKOUT3_GATE_EN                (1'b0),
//     .SC_CLKOUT4_GATE_EN                (1'b0),
//     .SC_CLKOUTPHY_GATE_EN              (1'b1),
//     .SC_CP_CUR_SEL                     (4'b0000),
//     .SC_CP_SELFBIAS_SEL                (2'b00),
//     .SC_DLDO_LOAD_CTRL                 (1'b0),
//     .SC_DLDO_TEST                      (2'b10),
//     .SC_DLDO_TEST_EN                   (1'b0),
//     .SC_DLDO_VREF_ADJ                  (3'b000),
//     .SC_DLDO_VREF_SEL                  (4'b0000),
//     .SC_DYNSEL_ENABLE                  (1'b0),
//     .SC_FDIV_CPHASE                    (7'd0),
//     .SC_FDIV_DUTY                      (FDIV),
//     .SC_FDIV_FPHASE                    (3'd0),
//     .SC_FDIV_MUXSEL_EN                 (1'b1),
//     .SC_FDIV_RATIO                     (FDIV),
//     .SC_FEEDBK_SEL                     (4'b0000),
//     .SC_FREQDETECT_BYPASSREXT_EN       (1'b0),
//     .SC_FREQDETECT_BYPASSR_EXT         (1'b0),
//     .SC_FREQDETECT_EN                  (1'b1),
//     .SC_FREQ_LOCKDET_MODE_SEL          (1'b0),
//     .SC_FREQ_LOCKDET_RSTNCTRL          (1'b0),
//     .SC_FREQ_LOCKDET_SET               (5'd28),
//     .SC_GLOGEN_ENABLE                  (1'b1),
//     .SC_ICP_BASE_SEL                   (2'b00),
//     .SC_IDIV_RATIO                     (IDIV),      // idiv /2
//     .SC_LDO_R_BYPASS_ENABLE            (1'b0),
//     .SC_LOCK_FILTER_PD                 (1'b1),
//     .SC_LPF_C                          (1'b0),
//     .SC_LPF_R                          (3'b000),
//     .SC_MDIV_RATIO                     (8'd1),
//     .SC_ODIV0_CPHASE                   (7'd0),
//     .SC_ODIV0_DUTY                     (ODIV0),
//     .SC_ODIV0_FPHASE                   (3'd0),
//     .SC_ODIV0_MUXSEL_EN                (1'b1),
//     .SC_ODIV0_RATIO                    (ODIV0),
//     .SC_ODIV1_CPHASE                   (7'd0),
//     .SC_ODIV1_DUTY                     (ODIV1),
//     .SC_ODIV1_FPHASE                   (3'd0),
//     .SC_ODIV1_MUXSEL_EN                (1'b1),
//     .SC_ODIV1_RATIO                    (ODIV1),
//     .SC_ODIV2_CPHASE                   (7'd0),
//     .SC_ODIV2_DUTY                     (ODIV2),
//     .SC_ODIV2_FPHASE                   (3'd0),
//     .SC_ODIV2_MUXSEL_EN                (1'b1),
//     .SC_ODIV2_RATIO                    (ODIV2),
//     .SC_ODIV3_CPHASE                   (7'd0),
//     .SC_ODIV3_DUTY                     (ODIV3),
//     .SC_ODIV3_FPHASE                   (3'd0),
//     .SC_ODIV3_MUXSEL_EN                (1'b1),
//     .SC_ODIV3_RATIO                    (ODIV3),
//     .SC_ODIV4_CPHASE                   (7'd0),
//     .SC_ODIV4_DUTY                     (ODIV4),
//     .SC_ODIV4_FPHASE                   (3'd0),
//     .SC_ODIV4_MUXSEL_EN                (1'b1),
//     .SC_ODIV4_RATIO                    (ODIV4),
//     .SC_ODIVPHY_CPHASE                 (7'd0),
//     .SC_ODIVPHY_DUTY                   (ODIVPHY),
//     .SC_ODIVPHY_FPHASE                 (3'd0),
//     .SC_ODIVPHY_MUXSEL_EN              (1'b1),
//     .SC_ODIVPHY_RATIO                  (ODIVPHY),
//     .SC_PFDEN_ENABLE                   (1'b1),
//     .SC_PFDTOP_CLKTEST_EN              (1'b0),
//     .SC_PFDTOP_CLKTEST_SEL             (1'b0),
//     .SC_PFDTOP_LSTEST_SEL              (3'b000),
//     .SC_PFD_DEADZONE                   (2'b00),
//     .SC_PLL_PWD_ENABLE                 (1'b0),
//     .SC_PLL_RST_ENABLE                 (1'b1),       //pll_rst enable
//     .SC_PLL_USE_APB                    (1'b0),
//     .SC_PPLL_DCTEST_SEL                (2'b00),
//     .SC_PPLL_VCTRL_TEST_EN             (1'b0),
//     .SC_VCTRL_INIT                     (2'b00),   
//     .CLKFBOUT                          (),
//     .CLKFBOUTN                         (),
//     .CLKOUT0                           (clkout0),
//     .CLKOUT0N                          (clkout0n),
//     .CLKOUT1                           (),
//     .CLKOUT1N                          (),
//     .CLKOUT2                           (),
//     .CLKOUT2N                          (),
//     .CLKOUT3                           (),
//     .CLKOUT3N                          (),
//     .CLKOUT4                           (),
//     .CLKOUT4N                          (),
//     .CLKOUTPHY                         (clkoutphy),
//     .CLKOUTPHYN                        (clkoutphyn),
//     .DCTEST_OUT                        (),
//     .LDO_ANA_TEST_MUX                  (),
//     .LDO_DIG_TEST_MUX                  (),
//     .LOCKOUT_CAS                       (),
//     .PLL_LOCK                          (pll_lock),
//     .PPLL_VCTRL_TEST                   (),
//     .PRDATA                            (),
//     .PREADY                            (),
//     .TEST_SO                           (),
//     .PFDTOP_CLK_TEST                   (),
//     .PLL_LS_TEST                       (),
//     .VCC                               (VCC),
//     .VCCA_PPLL                         (VCC),
//     .VSS                               (VSS),
//     .VSSA_PPLL                         (VSS),
//     .CLKFBOUT_GATE                     (1'b0),
//     .CLKOUT0_GATE                      (1'b0),
//     .CLKOUT1_GATE                      (1'b0),
//     .CLKOUT2_GATE                      (1'b0),
//     .CLKOUT3_GATE                      (1'b0),
//     .CLKOUT4_GATE                      (1'b0),
//     .CLKOUTPHY_GATE                    (clkoutphy_gate),
//     .CLK_FB                            (1'b0),
//     .CLK_IN0                           (clk_in0),
//     .CLK_IN1                           (1'b0),
//     .DYNSEL_CLKIN                      (1'b0),
//     .GLOGEN                            (glogen),
//     .GRS_N                             (glogen),
//     .GWEN                              (1'b1),
//     .LOCKIN_CAS                        (1'b1),
//     .PADDR                             (5'd0),
//     .PCLK                              (1'b0),
//     .PENABLE                           (1'b0),
//     .PFDEN                             (1'b1),
//     .PLL_PWD                           (1'b0),
//     .PLL_RST                           (pll_rst),
//     .PORN_1P8                          (VCC),
//     .PRESETN                           (1'b0),
//     .PSEL                              (1'b0),
//     .PWDATA                            (16'd0),
//     .PWRITE                            (1'b0),
//     .TEST_CLK                          (1'b1),
//     .TEST_MODE_N                       (1'b1),
//     .TEST_RSTN                         (1'b1),
//     .TEST_SE_N                         (1'b1),
//     .TEST_SI                           (1'b1),
//     .VREF1_ALDO_PPLL                   (VCC),
//     .VREF1_DLDO_PPLL                   (VCC),
//     .VREF2_ALDO_PPLL                   (VCC),
//     .VREF2_DLDO_PPLL                   (VCC)
//   );


endmodule
