
`define CONTROLLER_PHY_MODE

`define AXI_STANDARD_EN

`define CS_N_EN
 
`define DQ0_EN
 
`define DQ1_EN

`define RAS_DQS_EN

`define WE_DQS_EN

`define BA0_DQS_EN

`define BA2_EN

`define A4_DQS_EN

`define A5_DQS_EN

`define A12_EN

`define A13_EN

`define A14_EN

`define DEVICE_100H_EN
