module npu_top_vcs#(
parameter INSN_WIDTH            = 128,
parameter AXI_S_AXI_BURSTLENGTH = 64,
parameter AXI_M_AXI_BURSTLENGTH = 64,
parameter AXI_OUTSTANDING_DEPTH = 8,
parameter AXI_M_AXI_ID_WIDTH    = 10,
parameter AXI_M_AXI_ADDR_WIDTH  = 64,
parameter AXI_M_AXI_USER_WIDTH  = 1,
parameter AXI_M_AXI_DATA_WIDTH  = 256,
parameter DATA_AXI_ID_WIDTH     = 10,
parameter INSN_AXI_ID_WIDTH     = 10,
parameter AXI_S_AXI_ADDR_WIDTH  = 64,
parameter AXI_S_AXI_USER_WIDTH  = 1,
parameter AXI_S_AXI_DATA_WIDTH  = 256,
parameter PERI_DATA_WIDTH    = 256,
parameter PERI_ADDR_WIDTH    = 38,
parameter PERI_BUSRSTS_WIDTH = 22,
parameter SRAM_ADDR_WIDTH    = 20,
parameter AXI_M_AXI_DATA_BYTES   = AXI_M_AXI_DATA_WIDTH / 8,
parameter AXI_S_AXI_ID_WIDTH     = 10,
parameter AXI_S_AXI_DATA_BYTES   = AXI_S_AXI_DATA_WIDTH / 8,
parameter IFMAP_DMA_WIDTH         = 256,
parameter WEIGHT_DMA_WIDTH        = 256,
parameter VCUPARA_DMA_WIDTH       = 512,
parameter VCURES_DMA_WIDTH        = 256,
parameter OFMAP_DMA_WIDTH         = 256,
parameter IFMAP_WIDTH             = 128,
parameter WEIGHT_WIDTH            = 128,
parameter PSUM_WIDTH              = 512,
parameter VCUCODE_WIDTH           = 64,
parameter VCUPARA_WIDTH           = 256,
parameter VCURES_WIDTH            = 128,
parameter OFMAP_WIDTH             = 128,
parameter IFMAP_ADDR_BITS         = 14,
parameter WEIGHT_ADDR_BITS        = 15,
parameter PSUM_ADDR_BITS          = 11,
parameter VCUCODE_ADDR_BITS       = 7,
parameter VCUPARA_ADDR_BITS       = 8,
parameter VCURES_ADDR_BITS        = 13,
parameter OFMAP_ADDR_BITS         = 13,
parameter SYNCHRONIZE_FIFO_DEPTH = 128,
parameter integer INSN_ADDR_WIDTH    = 64,
parameter integer INSN_BUSRSTS_WIDTH = 8,
parameter integer INSN_DATA_WIDTH    = 256,
parameter integer INSN_FIFO_DEPTH    = 108,
parameter REG_WIDTH                  = 32,
parameter REG_NUM_BITS               = 8,
parameter SYNCHRONIZE_INSNBITS    = 128
)(
input clk, axi_clk, axi_rst_n, rst_n,
input       [AXI_S_AXI_ID_WIDTH-1:0]   axi_S_AXI_ARID,
input       [AXI_S_AXI_ADDR_WIDTH-1:0] axi_S_AXI_ARADDR,
input       [7:0]                      axi_S_AXI_ARLEN,
input       [2:0]                      axi_S_AXI_ARSIZE,
input       [1:0]                      axi_S_AXI_ARBURST,
input                                  axi_S_AXI_ARLOCK,
input       [3:0]                      axi_S_AXI_ARCACHE,
input       [2:0]                      axi_S_AXI_ARPROT,
input       [3:0]                      axi_S_AXI_ARQOS,
input       [AXI_S_AXI_USER_WIDTH-1:0] axi_S_AXI_ARUSER,
input                                  axi_S_AXI_ARVALID,
output wire                            axi_S_AXI_ARREADY,
output wire [AXI_S_AXI_ID_WIDTH-1:0]   axi_S_AXI_RID,
output wire [AXI_S_AXI_DATA_WIDTH-1:0] axi_S_AXI_RDATA,
output wire [1:0]                      axi_S_AXI_RRESP,
output wire                            axi_S_AXI_RLAST,
output wire [AXI_S_AXI_USER_WIDTH-1:0] axi_S_AXI_RUSER,
output wire                            axi_S_AXI_RVALID,
input                                  axi_S_AXI_RREADY,
input       [AXI_S_AXI_ID_WIDTH-1:0]   axi_S_AXI_AWID,
input       [AXI_M_AXI_ADDR_WIDTH-1:0] axi_S_AXI_AWADDR,
input       [7:0]                      axi_S_AXI_AWLEN,
input       [2:0]                      axi_S_AXI_AWSIZE,
input       [1:0]                      axi_S_AXI_AWBURST,
input                                  axi_S_AXI_AWLOCK,
input       [3:0]                      axi_S_AXI_AWCACHE,
input       [2:0]                      axi_S_AXI_AWPROT,
input       [3:0]                      axi_S_AXI_AWQOS,
input       [AXI_S_AXI_USER_WIDTH-1:0] axi_S_AXI_AWUSER,
input                                  axi_S_AXI_AWVALID,
output wire                            axi_S_AXI_AWREADY,
input       [AXI_S_AXI_DATA_WIDTH-1:0] axi_S_AXI_WDATA,
input       [AXI_S_AXI_DATA_BYTES-1:0] axi_S_AXI_WSTRB,
input                                  axi_S_AXI_WLAST,
input       [AXI_S_AXI_USER_WIDTH-1:0] axi_S_AXI_WUSER,
input                                  axi_S_AXI_WVALID,
output wire                            axi_S_AXI_WREADY,
output wire [AXI_S_AXI_ID_WIDTH-1:0]   axi_S_AXI_BID,
output wire [1:0]                      axi_S_AXI_BRESP,
output wire [AXI_S_AXI_USER_WIDTH-1:0] axi_S_AXI_BUSER,
output wire                            axi_S_AXI_BVALID,
input                                  axi_S_AXI_BREADY,
output wire [DATA_AXI_ID_WIDTH-1:0]    data_M_AXI_AWID,
output wire [AXI_M_AXI_ADDR_WIDTH-1:0] data_M_AXI_AWADDR,
output wire [7:0]                      data_M_AXI_AWLEN,
output wire [2:0]                      data_M_AXI_AWSIZE,
output wire [1:0]                      data_M_AXI_AWBURST,
output wire                            data_M_AXI_AWLOCK,
output wire [3:0]                      data_M_AXI_AWCACHE,
output wire [2:0]                      data_M_AXI_AWPROT,
output wire [3:0]                      data_M_AXI_AWQOS,
output wire [AXI_M_AXI_USER_WIDTH-1:0] data_M_AXI_AWUSER,
output wire                            data_M_AXI_AWVALID,
input                                  data_M_AXI_AWREADY,
output wire [AXI_M_AXI_DATA_WIDTH-1:0] data_M_AXI_WDATA,
output wire [AXI_M_AXI_DATA_BYTES-1:0] data_M_AXI_WSTRB,
output wire                            data_M_AXI_WLAST,
output wire [AXI_M_AXI_USER_WIDTH-1:0] data_M_AXI_WUSER,
output wire                            data_M_AXI_WVALID,
input                                  data_M_AXI_WREADY,
input       [DATA_AXI_ID_WIDTH-1:0]    data_M_AXI_BID,
input       [1:0]                      data_M_AXI_BRESP,
input       [AXI_M_AXI_USER_WIDTH-1:0] data_M_AXI_BUSER,
input                                  data_M_AXI_BVALID,
output wire                            data_M_AXI_BREADY,
output wire [DATA_AXI_ID_WIDTH-1:0]    data_M_AXI_ARID,
output wire [AXI_M_AXI_ADDR_WIDTH-1:0] data_M_AXI_ARADDR,
output wire [7:0]                      data_M_AXI_ARLEN,
output wire [2:0]                      data_M_AXI_ARSIZE,
output wire [1:0]                      data_M_AXI_ARBURST,
output wire                            data_M_AXI_ARLOCK,
output wire [3:0]                      data_M_AXI_ARCACHE,
output wire [2:0]                      data_M_AXI_ARPROT,
output wire [3:0]                      data_M_AXI_ARQOS,
output wire [AXI_M_AXI_USER_WIDTH-1:0] data_M_AXI_ARUSER,
output wire                            data_M_AXI_ARVALID,
input                                  data_M_AXI_ARREADY,
input       [DATA_AXI_ID_WIDTH-1:0]    data_M_AXI_RID,
input       [AXI_M_AXI_DATA_WIDTH-1:0] data_M_AXI_RDATA,
input       [1:0]                      data_M_AXI_RRESP,
input                                  data_M_AXI_RLAST,
input       [AXI_M_AXI_USER_WIDTH-1:0] data_M_AXI_RUSER,
input                                  data_M_AXI_RVALID,
output wire                            data_M_AXI_RREADY,
output wire [INSN_AXI_ID_WIDTH-1:0]    insn_M_AXI_AWID,
output wire [AXI_M_AXI_ADDR_WIDTH-1:0] insn_M_AXI_AWADDR,
output wire [7:0]                      insn_M_AXI_AWLEN,
output wire [2:0]                      insn_M_AXI_AWSIZE,
output wire [1:0]                      insn_M_AXI_AWBURST,
output wire                            insn_M_AXI_AWLOCK,
output wire [3:0]                      insn_M_AXI_AWCACHE,
output wire [2:0]                      insn_M_AXI_AWPROT,
output wire [3:0]                      insn_M_AXI_AWQOS,
output wire [AXI_M_AXI_USER_WIDTH-1:0] insn_M_AXI_AWUSER,
output wire                            insn_M_AXI_AWVALID,
input                                  insn_M_AXI_AWREADY,
output wire [AXI_M_AXI_DATA_WIDTH-1:0] insn_M_AXI_WDATA,
output wire [AXI_M_AXI_DATA_BYTES-1:0] insn_M_AXI_WSTRB,
output wire                            insn_M_AXI_WLAST,
output wire [AXI_M_AXI_USER_WIDTH-1:0] insn_M_AXI_WUSER,
output wire                            insn_M_AXI_WVALID,
input                                  insn_M_AXI_WREADY,
input       [DATA_AXI_ID_WIDTH-1:0]    insn_M_AXI_BID,
input       [1:0]                      insn_M_AXI_BRESP,
input       [AXI_M_AXI_USER_WIDTH-1:0] insn_M_AXI_BUSER,
input                                  insn_M_AXI_BVALID,
output wire                            insn_M_AXI_BREADY,
output wire [INSN_AXI_ID_WIDTH-1:0]    insn_M_AXI_ARID,
output wire [AXI_M_AXI_ADDR_WIDTH-1:0] insn_M_AXI_ARADDR,
output wire [7:0]                      insn_M_AXI_ARLEN,
output wire [2:0]                      insn_M_AXI_ARSIZE,
output wire [1:0]                      insn_M_AXI_ARBURST,
output wire                            insn_M_AXI_ARLOCK,
output wire [3:0]                      insn_M_AXI_ARCACHE,
output wire [2:0]                      insn_M_AXI_ARPROT,
output wire [3:0]                      insn_M_AXI_ARQOS,
output wire [AXI_M_AXI_USER_WIDTH-1:0] insn_M_AXI_ARUSER,
output wire                            insn_M_AXI_ARVALID,
input                                  insn_M_AXI_ARREADY,
input       [INSN_AXI_ID_WIDTH-1:0]    insn_M_AXI_RID,
input       [AXI_M_AXI_DATA_WIDTH-1:0] insn_M_AXI_RDATA,
input       [1:0]                      insn_M_AXI_RRESP,
input                                  insn_M_AXI_RLAST,
input       [AXI_M_AXI_USER_WIDTH-1:0] insn_M_AXI_RUSER,
input                                  insn_M_AXI_RVALID,
output wire                            insn_M_AXI_RREADY
);
endmodule